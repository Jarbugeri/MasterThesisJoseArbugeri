LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY PROTECAO IS
	PORT (
		CLK : IN STD_LOGIC;
		RESET : IN STD_LOGIC;
		PWMAin : IN STD_LOGIC;
		PWMBin : IN STD_LOGIC;
		OverC : IN STD_LOGIC;
		CORRENTE_mA : IN SIGNED (23 DOWNTO 0);
		TENSAO_mV : IN UNSIGNED (23 DOWNTO 0);
		CORRENTE_MAX : OUT SIGNED (23 DOWNTO 0);
		OVERTENSION : OUT STD_LOGIC;
		OverC_HARDWARE : OUT STD_LOGIC;
		OverC_SOFTWARE : OUT STD_LOGIC;
		ENABLEP : OUT STD_LOGIC;
		ENABLEN : OUT STD_LOGIC;
		PWMPout : OUT STD_LOGIC;
		PWMNout : OUT STD_LOGIC);
END PROTECAO;

ARCHITECTURE ARCH OF PROTECAO IS

	--REGISTER
	SIGNAL FLAG_CORRENTE : STD_LOGIC := '0';
	SIGNAL FLAG_TENSAO : STD_LOGIC := '0';
	SIGNAL FLAG_OVERC : STD_LOGIC := '0';
	CONSTANT LIMITE_CORRENTE_P : SIGNED (23 DOWNTO 0) := TO_SIGNED( 15000, 24); --vALOR EM mA 
	CONSTANT LIMITE_CORRENTE_N : SIGNED (23 DOWNTO 0) := TO_SIGNED(-15000, 24); --vALOR EM mA 
	CONSTANT LIMITE_TENSAO : UNSIGNED (23 DOWNTO 0) := TO_UNSIGNED(200000, 24); --vALOR EM mV 
	SIGNAL CORRENTE_VALUE : SIGNED (23 DOWNTO 0) := TO_SIGNED( 0, 24);

BEGIN

	OVERTENSION <= FLAG_TENSAO;
	OverC_HARDWARE <= FLAG_OVERC;
	OverC_SOFTWARE <= FLAG_CORRENTE;
	CORRENTE_MAX <= CORRENTE_VALUE;

	PROCESS (CLK, RESET) BEGIN
		IF (RESET = '1') THEN
			FLAG_CORRENTE <= '0';
			FLAG_TENSAO <= '0';
			FLAG_OVERC <= '0';
			PWMPout <= '0';
			PWMNout <= '0';
			ENABLEP <= '0';
			ENABLEN <= '0';
			CORRENTE_VALUE <= TO_SIGNED( 0, 24);
		ELSIF RISING_EDGE(CLK) THEN

			IF CORRENTE_mA > LIMITE_CORRENTE_P THEN
				FLAG_CORRENTE <= '1';
				CORRENTE_VALUE <= CORRENTE_mA;
			END IF;

			IF CORRENTE_mA < LIMITE_CORRENTE_N THEN
				FLAG_CORRENTE <= '1';
				CORRENTE_VALUE <= CORRENTE_mA;
			END IF;

			IF TENSAO_mV >= LIMITE_TENSAO THEN
				FLAG_TENSAO <= '1';
			END IF;

			IF OverC = '0' THEN -- OverC == 1, Iin < 20 A , OverC == 0, Iin > 20 A
				FLAG_OVERC <= '1';
			END IF;

			IF FLAG_CORRENTE = '1' OR FLAG_TENSAO = '1' THEN -- OR FLAG_OVERC = '1' Removi pq ta com ruido
				PWMPout <= '0';
				PWMNout <= '0';
				ENABLEP <= '0';
				ENABLEN <= '0';
			ELSE
				PWMPout <= PWMAin;
				PWMNout <= PWMBin;
				ENABLEP <= '1';
				ENABLEN <= '1';
			END IF;
		END IF;
	END PROCESS;
END ARCH;